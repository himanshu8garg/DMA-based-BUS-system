library IEEE;
  use IEEE.std_logic_1164.all;
  use work.ensc350_package.all;
  use ieee.numeric_std.all;
  
entity ensc350 is
  port(  	clk,resetn           : in  Std_logic;
			iaddr_out            : out Std_logic_vector(iaddr_size-1 downto 0);
			idata_in             : in  Std_logic_vector(instr_size-1 downto 0);
			daddr_out            : out Std_logic_vector(daddr_size-1 downto 0);
			dmem_read,dmem_write : out std_logic;
			ddata_in             : in  Std_logic_vector(data_size-1  downto 0);
			ddata_out            : out Std_logic_vector(data_size-1  downto 0));
end ensc350;

architecture struct of ensc350 is

component rfile
	generic( size      : positive := 32; addr_size : positive := 5 );  
	port(  clk,resetn   : in  Std_logic;
           ra,rb        : in  Std_logic_vector(addr_size-1 downto 0);
           a_out,b_out  : out Std_logic_vector(size-1 downto 0);
           rd1          : in  Std_logic_vector(addr_size-1 downto 0);
           d1_in        : in  Std_logic_vector(size-1 downto 0) ); 
end component;

component full_alu
    generic (size : integer := 16);
    port(  in1,in2       : in  std_logic_vector(size-1 downto 0);
           op            : in  alu_commands;
           result        : out Std_logic_vector(size-1 downto 0);
           overflow      : out Std_logic );
end component;

component mem_control
  port ( -- Communication to the processor: Operation to be performed, Data to be stored, data read
         mem_op                : in  mem_commands;
		 addr_base,addr_offset : in  std_logic_vector(data_size-1 downto 0);
		 store_data    		   : in  std_logic_vector(data_size-1 downto 0);
         read_data     		   : out std_logic_vector(data_size-1 downto 0);
		 -- Bus control: Output address, Control Signals, Data Out and Data In (Note: Signals with capital letters 
		 -- connect out of the  processor. Note: On-Chip Bus CAN NEVER BE BIDIRECTIONAL, has to be either IN or OUT
         ADDR_OUT      : out std_logic_vector(daddr_size-1 downto 0);
		 MR, MW        : out std_logic;
         DATA_IN       : in  std_logic_vector(data_size-1 downto 0);
         DATA_OUT      : out std_logic_vector(data_size-1 downto 0)  );   
end component;

component decodeop
    port( instr                        : in   Std_logic_vector(instr_size-1 downto 0);
          rs1,rs2,rd                   : out  Std_logic_vector(rf_addr_size-1 downto 0);
          pc_op                        : out  pc_commands;
          alu_op                       : out  alu_commands;
          mul_op                       : out  mul_commands;
		  mem_op                       : out  mem_commands;
		  operand_sel                  : out  operand_select; 
          wb_sel                       : out  wb_select;
		  immediate                    : out  Std_logic_vector(data_size-1 downto 0);
          illegal_opcode               : out  Std_logic );
end component;

component pc_calc 
  port ( clk,resetn           : in  std_logic;
         pc_op                : in  pc_commands;
		 rs1,rs2              : in  std_logic_vector(data_size-1 downto 0);
		 offset               : in  std_logic_vector(data_size-1 downto 0);
		 IADDR_OUT            : out std_logic_vector(iaddr_size-1 downto 0) );   
end component;

component multiplier
  generic(size : positive :=16);
  port (in1,in2 : in  std_logic_vector(size-1 downto 0); 
        result  : out std_logic_vector(size-1 downto 0));
end component;

signal instr       : std_logic_vector(instr_size-1 downto 0);
signal rs1,rs2,rd1 : std_logic_vector(rf_addr_size-1 downto 0);
signal rf_out1,rf_out2,rf_in1,immediate,alu_in1,alu_in2,alu_out1,mem_out1,mul_out1 : std_logic_vector(data_size-1 downto 0);
signal alu_op      : alu_commands;
signal mul_op      : mul_commands; 
signal mem_op      : mem_commands;
signal pc_op       : pc_commands;
signal operand_sel : operand_select; 
signal wb_sel      : wb_select; 
signal exc_overflow, exc_illegal_opcode : std_logic;

--pipeline signals
signal Pipe_RD : std_logic_vector(3 downto 0);
signal Pipe_mul_out : std_logic_vector(data_size-1 downto 0);
signal Pipe_alu_out : std_logic_vector(data_size-1 downto 0);
signal Pipe_wb_sel : wb_select;
 
signal Pipe_instr : std_logic_vector(instr_size-1 downto 0);

begin

	intr_fetch : instr <= idata_in;
	
	-- Decodeop Logic
	instr_decode : decodeop port map (instr,rs1,rs2,rd1,
	                                  pc_op,alu_op,mul_op,mem_op,
									  operand_sel,wb_sel,immediate,exc_illegal_opcode);
									  
	pc_calculation : pc_calc port map (clk,resetn,pc_op,rf_out1,rf_out2,immediate,
	                                   IADDR_OUT); 


    -- Register File: 32-slots of 16 bits, r0 is always zero
	register_file : rfile generic map (size=>data_size, addr_size=>rf_addr_size)
	                      port map (clk,resetn,rs1,rs2,rf_out1,rf_out2,
									Pipe_RD,rf_in1);
									
	-- Alu Operand Selection								
	alu_in2_mux : alu_in2 <= immediate when operand_sel=operand_immed else rf_out2;
	alu_in1_mux : alu_in1 <= rf_out1;
	
	-- Alu: Includes shifting operations							
	alu1 : full_alu generic map (size=>data_size)
	                port map (alu_in1,alu_in2,alu_op,alu_out1,exc_overflow);
					
	-- Multiplier: 
     mult : multiplier generic map (size=>data_size)
	                   port map (rf_out1,rf_out2,mul_out1);
	 
	-- Memory Control Logic
	memory_logic : mem_control port map (mem_op,rf_out1,immediate,rf_out2,mem_out1,
	                                     DADDR_OUT,DMEM_READ,DMEM_WRITE,DDATA_IN,DDATA_OUT);
 
	wb_mux : rf_in1 <= Pipe_alu_out when Pipe_wb_sel=wb_alu else 
	                   ddata_in when Pipe_wb_sel=wb_mem else
			   Pipe_mul_out when Pipe_wb_sel=wb_mul else				
			   (others=>'0');

	pipeline: process(clk,resetn)
	begin
		if resetn = '0' then
			Pipe_RD<=x"0";
			Pipe_mul_out<=x"00000000";
			Pipe_alu_out<=x"00000000";
			Pipe_wb_sel<=wb_alu;
			Pipe_instr<=x"00000000";
		else if clk'event and clk='1' then 
	 		Pipe_RD<=rd1;
			Pipe_mul_out<=mul_out1;
			Pipe_alu_out<=alu_out1;
			Pipe_wb_sel<=wb_sel;
			Pipe_instr<=instr;
		end if; 
	end if;

	end process;	
end struct;